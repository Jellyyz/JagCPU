module mem_wb #(parameter width = 32)
(
    input clk,
    input rst

);

endmodule : mem_wb 