import rv32i_types::*;

module EX(

); 


endmodule 
