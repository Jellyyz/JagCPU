module ex_mem #(parameter width = 32)
(
    input clk,
    input rst

);

endmodule : ex_mem 