module branch_predictor (

    input clk, rst


    



); 




endmodule  

