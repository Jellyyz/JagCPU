import rv32i_types::*;

module EX_MEM(

); 


endmodule 
