module cache(



); 


endmodule 